`timescale 1ns / 1ps

module pipeline (
					input wire clk,
					input wire rst_n
				);
