`timescale 1ns /1ps

module instruction_fetch(
						input wire 	clk,
						input wire 	rst_n,
						input wire
					
